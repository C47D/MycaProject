library verilog;
use verilog.vl_types.all;
entity mrm is
    port(
        a               : in     vl_logic_vector(3 downto 0);
        D               : out    vl_logic_vector(6 downto 0)
    );
end mrm;
