library verilog;
use verilog.vl_types.all;
entity MycaII_vlg_vec_tst is
end MycaII_vlg_vec_tst;
