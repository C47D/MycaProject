library verilog;
use verilog.vl_types.all;
entity um1b_vlg_vec_tst is
end um1b_vlg_vec_tst;
