library verilog;
use verilog.vl_types.all;
entity myca1_vlg_vec_tst is
end myca1_vlg_vec_tst;
