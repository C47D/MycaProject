library verilog;
use verilog.vl_types.all;
entity usomycaII_vlg_vec_tst is
end usomycaII_vlg_vec_tst;
