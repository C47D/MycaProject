library verilog;
use verilog.vl_types.all;
entity div_vlg_check_tst is
    port(
        ck1s            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end div_vlg_check_tst;
