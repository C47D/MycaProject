library verilog;
use verilog.vl_types.all;
entity mrm_vlg_vec_tst is
end mrm_vlg_vec_tst;
