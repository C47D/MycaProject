library verilog;
use verilog.vl_types.all;
entity um1bb_vlg_vec_tst is
end um1bb_vlg_vec_tst;
