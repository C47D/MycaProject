library verilog;
use verilog.vl_types.all;
entity sumador_vlg_sample_tst is
    port(
        ci              : in     vl_logic;
        pc              : in     vl_logic_vector(7 downto 0);
        sampler_tx      : out    vl_logic
    );
end sumador_vlg_sample_tst;
