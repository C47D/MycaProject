library verilog;
use verilog.vl_types.all;
entity div_vlg_sample_tst is
    port(
        ck              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end div_vlg_sample_tst;
