library verilog;
use verilog.vl_types.all;
entity dr_vlg_vec_tst is
end dr_vlg_vec_tst;
